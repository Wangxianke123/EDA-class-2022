TestBench2 for Homework3 

Vin 1 0 3
R1 1 2 2k
R2 2 0 100
C1 2 0 2e-10

.DC Vin 0.5 2 0.1
.Print DC V(2)
.end
