TestBench3 for Homework4
* 2022-10-17
* Origin: Lecture 6 Circuit III Page-14

R1 1 0 5
G2 1 0 1 2 2
R3 1 2 6
R4 2 0 8
Is 0 2 10
Vs 3 2 1
R8 3 4 5
E7 4 0 1 2 13
.DC VS 1 2 0.1
.END
