TestBench1 for Homework3 
* 2022 EDA course testbench netlist  
Vin 1 0 3
R1 1 2 200
R2 2 0 100
.op
.end